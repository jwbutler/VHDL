-- THIS MAY COMPILE, BUT I'M NOT SURE IT DOES ANYTHING.
-- ADD MORE STUFFS TO IT
-- MAYBE MAKE SOME SCHEMATICS (FIRST)?

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE WORK.ALL;

ENTITY PROCESSOR IS
	PORT(CLK: IN STD_LOGIC;
			 DIN: IN STD_LOGIC_VECTOR (0 TO 15);
			 RUN: IN STD_LOGIC;
			 RESET: IN STD_LOGIC;
			 U_BUS: INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
			 DONE: OUT STD_LOGIC);
END PROCESSOR;

ARCHITECTURE BEHV OF PROCESSOR IS
	COMPONENT REGISTER_9
		PORT (CLK: IN STD_LOGIC;
					EN: IN STD_LOGIC;
					D: IN STD_LOGIC_VECTOR(0 TO 8);
					Q: OUT STD_LOGIC_VECTOR(0 TO 8));
	END COMPONENT;
	COMPONENT REGISTER_16
		PORT (CLK: IN STD_LOGIC;
  	  	  EN: IN STD_LOGIC;
    	    D: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
     		  Q: OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
	END COMPONENT;
	COMPONENT ADDER
		PORT (X: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
 					Y: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
					Z: OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
	END COMPONENT;
	COMPONENT SUB
		PORT (X: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
					Y: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
					Z: OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
	END COMPONENT;
	COMPONENT COUNTER
		PORT (CLR: IN STD_LOGIC;
					CLK: IN STD_LOGIC;
					Q: INOUT STD_LOGIC_VECTOR (0 TO 1));
	END COMPONENT;
	COMPONENT CONTROL
		PORT(RUN: IN STD_LOGIC;
				 RESETN: IN STD_LOGIC;
				 INS: IN STD_LOGIC_VECTOR(0 TO 8); -- TO OR DOWNTO?
				 CNT: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
				 A_IN: OUT STD_LOGIC;
				 CLR: OUT STD_LOGIC;
				 DONE: OUT STD_LOGIC;
				 DIN_OUT: OUT STD_LOGIC;
				 G_IN: OUT STD_LOGIC;
				 G_OUT: OUT STD_LOGIC;
				 IR_IN: OUT STD_LOGIC;
				 R_IN: OUT STD_LOGIC_VECTOR(0 TO 7); -- TO OR DOWNTO?
				 R_OUT: OUT STD_LOGIC_VECTOR(0 TO 7);
				 ADDSUB: OUT STD_LOGIC); -- TO OR DOWNTO?
	END COMPONENT;
	COMPONENT MUX10TO1
     PORT(
       RN: IN STD_LOGIC_VECTOR(0 TO 7);
       I0: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
       I1: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
       I2: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
       I3: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
       I4: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
       I5: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
       I6: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
       I7: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
       DIN: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
       G: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
       D: IN STD_LOGIC;
       GOUT: IN STD_LOGIC;
  		 O: OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
     );
	END COMPONENT;
	COMPONENT ADDSUB
		PORT (X, Y: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
			SUB: IN STD_LOGIC; -- 1 = subtract mode
			F: OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
	END COMPONENT;
	SIGNAL CLR: STD_LOGIC;
	SIGNAL A_IN: STD_LOGIC;
	SIGNAL DIN_OUT: STD_LOGIC;
	SIGNAL G_IN: STD_LOGIC;
	SIGNAL G_OUT: STD_LOGIC;
	SIGNAL IR_IN: STD_LOGIC;
	SIGNAL EN_ADDSUB: STD_LOGIC;
	SIGNAL T: STD_LOGIC_VECTOR (0 TO 1);
	SIGNAL R_OUT: STD_LOGIC_VECTOR (0 TO 7);
	SIGNAL R_IN: STD_LOGIC_VECTOR (0 TO 7);
	SIGNAL R_DATA_OUT_0: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL R_DATA_OUT_1: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL R_DATA_OUT_2: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL R_DATA_OUT_3: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL R_DATA_OUT_4: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL R_DATA_OUT_5: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL R_DATA_OUT_6: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL R_DATA_OUT_7: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL INS: STD_LOGIC_VECTOR (0 TO 8);
	SIGNAL IR_OUT: STD_LOGIC_VECTOR (0 TO 8);
	SIGNAL A_OUT: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL G_OUT_DATA: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL ADDSUB_OUT: STD_LOGIC_VECTOR (15 DOWNTO 0);
BEGIN
	-- WHAT DOES THE U STAND FOR, ANYWAY
	U_COUNTER: COUNTER PORT MAP (CLR, CLK, T);
	U_CONTROL: CONTROL PORT MAP (RUN, RESET, INS, T, A_IN, CLR, DONE,
    DIN_OUT, G_IN, G_OUT, IR_IN, R_IN, R_OUT, EN_ADDSUB);

	U_IR: REGISTER_9 PORT MAP (CLK, IR_IN, INS, IR_OUT);
	U_A: REGISTER_16 PORT MAP (CLK, A_IN, U_BUS, A_OUT);
	U_G: REGISTER_16 PORT MAP (CLK, G_IN, ADDSUB_OUT, G_OUT_DATA);
	U_R0: REGISTER_16 PORT MAP (CLK, R_IN(0), U_BUS, R_DATA_OUT_0);
	U_R1: REGISTER_16 PORT MAP (CLK, R_IN(1), U_BUS, R_DATA_OUT_1);
	U_R2: REGISTER_16 PORT MAP (CLK, R_IN(2), U_BUS, R_DATA_OUT_2);
	U_R3: REGISTER_16 PORT MAP (CLK, R_IN(3), U_BUS, R_DATA_OUT_3);
	U_R4: REGISTER_16 PORT MAP (CLK, R_IN(4), U_BUS, R_DATA_OUT_4);
	U_R5: REGISTER_16 PORT MAP (CLK, R_IN(5), U_BUS, R_DATA_OUT_5);
	U_R6: REGISTER_16 PORT MAP (CLK, R_IN(6), U_BUS, R_DATA_OUT_6);
	U_R7: REGISTER_16 PORT MAP (CLK, R_IN(7), U_BUS, R_DATA_OUT_7);

	U_MUX: MUX10TO1 PORT MAP (R_OUT, R_DATA_OUT_0, R_DATA_OUT_1, R_DATA_OUT_2,
													R_DATA_OUT_3, R_DATA_OUT_4, R_DATA_OUT_5,
													R_DATA_OUT_6, R_DATA_OUT_7, DIN, G_OUT_DATA,
													DIN_OUT, G_OUT,	U_BUS);
	U_ADDSUB: ADDSUB PORT MAP (A_OUT, U_BUS, EN_ADDSUB, ADDSUB_OUT);
	
	PROCESS (DIN, CLK)
	BEGIN
		IF T="00" THEN
			INS(0) <= DIN(0);
			INS(1) <= DIN(1);
			INS(2) <= DIN(2);
			INS(3) <= DIN(3);
			INS(4) <= DIN(4);
			INS(5) <= DIN(5);
			INS(6) <= DIN(6);
			INS(7) <= DIN(7);
			INS(8) <= DIN(8);
		END IF;
	END PROCESS;
END BEHV;