LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY MUX10TO1 IS
     PORT(
       -- PARTY.
       RN: in STD_LOGIC_VECTOR(0 TO 7);
       I0: in STD_LOGIC_VECTOR(15 DOWNTO 0);
       I1: in STD_LOGIC_VECTOR(15 DOWNTO 0);
       I2: in STD_LOGIC_VECTOR(15 DOWNTO 0);
       I3: in STD_LOGIC_VECTOR(15 DOWNTO 0);
       I4: in STD_LOGIC_VECTOR(15 DOWNTO 0);
       I5: in STD_LOGIC_VECTOR(15 DOWNTO 0);
       I6: in STD_LOGIC_VECTOR(15 DOWNTO 0);
       I7: in STD_LOGIC_VECTOR(15 DOWNTO 0);
       DIN: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
       G: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
       D: IN STD_LOGIC;
       GOUT: IN STD_LOGIC;
       O: out STD_LOGIC_VECTOR(15 DOWNTO 0)
     );
   END  MUX10TO1;            
--architecture definition
   architecture behv of mux10to1 is
-- start of design
      SIGNAL ENABLES: STD_LOGIC_VECTOR(0 TO 9);
begin
  -- THIS PROCESS LOOPS THROUGH TO CONSTRUCT THE ENABLE 
	PROCESS (RN, I0, I1, I2, I3, I4, I5, I6, I7,DIN, G,D, GOUT)
	 BEGIN
	  FOR I IN 0 TO 7 LOOP
		  ENABLES(I) <= RN(I);
		END LOOP;
		ENABLES(8) <= D;
		ENABLES(9) <= GOUT;
	END PROCESS;
	-- FROM ENABLES CHOOSE WHICH OF THE INPUTS TO OUTPUT
	  WITH ENABLES  SELECT
		O <=      I0 WHEN "1000000000",
				  I1 WHEN "0100000000",
				  I2 WHEN "0010000000",
				  I3 WHEN "0001000000",
				  I4 WHEN "0000100000",
				  I5 WHEN "0000010000",
				  I6 WHEN "0000001000",
				  I7 WHEN "0000000100",
				  DIN WHEN "0000000010",
				  G WHEN "0000000001",
				  "XXXXXXXXXXXXXXXX" WHEN OTHERS;
end behv;
