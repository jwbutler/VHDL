LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE WORK.ALL;
--ENTITY DECLARATION
   ENTITY TESTMUX IS
   END TESTMUX;
--ARCHITECTURE DEFINITION
   ARCHITECTURE TB OF TESTMUX IS
--COMPONENT DECLARATION
   COMPONENT MUX10TO1 IS
   PORT( 		
	   -- PARTY.
		   RN: IN STD_LOGIC_VECTOR(0 TO 7);
		   I0: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		   I1: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		   I2: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		   I3: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		   I4: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		   I5: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		   I6: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		   I7: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		   DIN: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		   G: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		   D: IN STD_LOGIC;
		   GOUT: IN STD_LOGIC;
		   O: OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
        );
   END COMPONENT;
--SIGNAL DECLARATION
		   SIGNAL T_RN: STD_LOGIC_VECTOR(0 TO 7);
		   SIGNAL T_I0: STD_LOGIC_VECTOR(15 DOWNTO 0);
		   SIGNAL T_I1: STD_LOGIC_VECTOR(15 DOWNTO 0);
		   SIGNAL T_I2: STD_LOGIC_VECTOR(15 DOWNTO 0);
		   SIGNAL T_I3: STD_LOGIC_VECTOR(15 DOWNTO 0);
		   SIGNAL T_I4: STD_LOGIC_VECTOR(15 DOWNTO 0);
		   SIGNAL T_I5: STD_LOGIC_VECTOR(15 DOWNTO 0);
		   SIGNAL T_I6: STD_LOGIC_VECTOR(15 DOWNTO 0);
		   SIGNAL T_I7: STD_LOGIC_VECTOR(15 DOWNTO 0);
		   SIGNAL T_DIN: STD_LOGIC_VECTOR(15 DOWNTO 0);
		   SIGNAL T_G: STD_LOGIC_VECTOR(15 DOWNTO 0);
		   SIGNAL T_D: STD_LOGIC;
		   SIGNAL T_GOUT: STD_LOGIC;
		   SIGNAL T_O: STD_LOGIC_VECTOR(15 DOWNTO 0);
  BEGIN
    
--COMPONENT STATEMENTS (CONCURRENT STATEMENT )
      TESTMUX: MUX10TO1 PORT MAP (T_RN,T_I0,T_I1,T_I2,T_I3,T_I4,T_I5,T_I6,T_I7,T_DIN,T_G,T_D,T_GOUT,T_O); 
--PROCESS STATEMENTS
      PROCESS
--VARIABLE DECLARATION
      VARIABLE ERR_CNT: INTEGER := 0;
   BEGIN
     REPORT "STARTING!";
-- SETTING THE REGISTERS
	T_I0 <= "0101010101010101";
	T_I1 <= "0001110001110101";
	T_I2 <= "1110101010101010";
	T_I3 <= "1010101000011001";
	T_I4 <= "0000000000000000";
	T_I5 <= "1111111111111111";
	T_I6 <= "0000001000101010";
	T_I7 <= "1001001000100010";
	T_DIN <= "1000100100100001";
	T_G <= "1111111011110011";
	
--THE TEST CASE I0
  REPORT "STARTING!";
	T_RN <= "10000000";
	T_D <= '0';
	T_GOUT <= '0' ;
   WAIT FOR 2 NS;
   ASSERT (T_O = "0101010101010101") REPORT "I0 CASE IS INCORRECT!" SEVERITY ERROR;
   IF (T_O /= "0101010101010101") THEN
       ERR_CNT := ERR_CNT + 1;
   END IF;
   WAIT FOR 10 NS;
 
 --THE TEST CASE I1
	T_RN <= "01000000";
	T_D <= '0';
	T_GOUT <= '0';
   WAIT FOR 2 NS;
   ASSERT (T_O = "0001110001110101") REPORT "I1 CASE IS INCORRECT!" SEVERITY ERROR;
   IF (T_O /= "0001110001110101") THEN
       ERR_CNT := ERR_CNT + 1;
   END IF;
   WAIT FOR 10 NS;
   
 --THE TEST CASE I2
	T_RN <= "00100000";
	T_D <= '0';
	T_GOUT <= '0';
   WAIT FOR 2 NS;
   ASSERT (T_O = "1110101010101010") REPORT "I2 CASE IS INCORRECT!" SEVERITY ERROR;
   IF (T_O /= "1110101010101010") THEN
       ERR_CNT := ERR_CNT + 1;
   END IF;
   WAIT FOR 10 NS;

 --THE TEST CASE I3
	T_RN <= "00010000";
	T_D <= '0';
	T_GOUT <= '0';
   WAIT FOR 2 NS;
   ASSERT (T_O = "1010101000011001") REPORT "I3 CASE IS INCORRECT!" SEVERITY ERROR;
   IF (T_O /= "1010101000011001") THEN
       ERR_CNT := ERR_CNT + 1;
   END IF;
   WAIT FOR 10 NS;
   
  --THE TEST CASE I4
	T_RN <= "00001000";
	T_D <= '0';
	T_GOUT <= '0';
   WAIT FOR 2 NS;
   ASSERT (T_O = "0000000000000000") REPORT "I4 CASE IS INCORRECT!" SEVERITY ERROR;
   IF (T_O /= "0000000000000000") THEN
       ERR_CNT := ERR_CNT + 1;
   END IF;
   WAIT FOR 10 NS;
   
   --THE TEST CASE I5
	T_RN <= "00000100";
	T_D <= '0';
	T_GOUT <= '0' ;
   WAIT FOR 2 NS;
   ASSERT (T_O = "1111111111111111") REPORT "I5 CASE IS INCORRECT!" SEVERITY ERROR;
   IF (T_O /= "1111111111111111") THEN
       ERR_CNT := ERR_CNT + 1;
   END IF;
   WAIT FOR 10 NS;  
 
    --THE TEST CASE I6
	T_RN <= "00000010";
	T_D <= '0';
	T_GOUT <= '0' ;
   WAIT FOR 2 NS;
   ASSERT (T_O = "0000001000101010") REPORT "I6 CASE IS INCORRECT!" SEVERITY ERROR;
   IF (T_O /= "0000001000101010") THEN
       ERR_CNT := ERR_CNT + 1;
   END IF;
   WAIT FOR 10 NS;

    --THE TEST CASE I7
	T_RN <= "00000001";
	T_D <= '0';
	T_GOUT <= '0' ;
   WAIT FOR 2 NS;
   ASSERT (T_O = "1001001000100010") REPORT "I7 CASE IS INCORRECT!" SEVERITY ERROR;
   IF (T_O /= "1001001000100010") THEN
       ERR_CNT := ERR_CNT + 1;
   END IF;
   WAIT FOR 10 NS;

    --THE TEST CASE D
	T_RN <= "00000000";
	T_D <= '1';
	T_GOUT <= '0' ;
   WAIT FOR 2 NS;
   ASSERT (T_O = "1000100100100001") REPORT "D CASE IS INCORRECT!" SEVERITY ERROR;
   IF (T_O /= "1000100100100001") THEN
       ERR_CNT := ERR_CNT + 1;
   END IF;
   WAIT FOR 10 NS;

    --THE TEST CASE GOUT
	T_RN <= "00000000";
	T_D <= '0';
	T_GOUT <= '1' ;
   WAIT FOR 2 NS;
   ASSERT (T_O = "1111111011110011") REPORT "GOUT CASE IS INCORRECT!" SEVERITY ERROR;
   IF (T_O /= "1111111011110011") THEN
       ERR_CNT := ERR_CNT + 1;
   END IF;
   WAIT FOR 10 NS;   
   
-- SUMMARY OF ALL THE TEST CASES
-- 	REPORT "SUMMARY!";
   IF (ERR_CNT=0) THEN
      ASSERT FALSE
      REPORT "TESTBENCH OF MUX10TO1 COMPLETED SUCCESSFULLY!"
      SEVERITY NOTE;
   ELSE
      ASSERT FALSE
      REPORT "SOMETHING WRONG, TRY TEST AGAIN"
      SEVERITY ERROR;
   END IF;
   WAIT;
 END PROCESS;
END TB;
--CONFIGURATION DECLARATION
CONFIGURATION CFG_TB OF TESTMUX IS
FOR TB
END FOR;
END CFG_TB;
