LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ADDSUB IS
	PORT (X: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
				Y: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
				SUB: IN STD_LOGIC; -- 1 = subtract mode
				F: OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
END ADDSUB;

ARCHITECTURE BEHV OF ADDSUB IS
	COMPONENT ADDER
		PORT (X: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
					Y: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
					Z: OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
	END COMPONENT;
	COMPONENT SUBTRACTOR
		PORT (X: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
					Y: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
					Z: OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
	END COMPONENT;
	SIGNAL Z_ADD: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL Z_SUB: STD_LOGIC_VECTOR (15 DOWNTO 0);
BEGIN
	U_ADDER: ADDER PORT MAP (X, Y, Z_ADD);
	U_SUB: SUBTRACTOR PORT MAP (X, Y, Z_SUB);
	
	PROCESS (X, Y, SUB, Z_ADD, Z_SUB)
	BEGIN
		IF SUB='0' THEN
			F <= Z_ADD;
		ELSE
			F <= Z_SUB;
		END IF;
	END PROCESS;
END BEHV;