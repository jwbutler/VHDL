LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY REGISTER_9 IS
	PORT (CLK: IN STD_LOGIC;
				EN: IN STD_LOGIC;
				D: IN STD_LOGIC_VECTOR(0 TO 8);
				Q: OUT STD_LOGIC_VECTOR(0 TO 8));
END REGISTER_9;

ARCHITECTURE BEHV OF REGISTER_9 IS
BEGIN
	PROCESS (D, EN, CLK)
	BEGIN
    IF EN='1' AND CLK' EVENT AND (NOT (NOT CLK))='1' THEN
			Q <= D;
    END IF;
	END PROCESS;
END BEHV;