LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY T_FF IS
	PORT (EN: IN STD_LOGIC;
				T: IN STD_LOGIC;
				Q: INOUT STD_LOGIC := '0');
END T_FF;

ARCHITECTURE BEHV OF T_FF IS
BEGIN
	PROCESS(EN, T)
	BEGIN
		IF EN='1' AND T='1' AND T' EVENT THEN
			Q <= NOT Q;
		END IF;
	END PROCESS;
END BEHV;