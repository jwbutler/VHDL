LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DECODER_3_8 IS
	PORT (I: IN STD_LOGIC_VECTOR(2 DOWNTO 0);	-- TO OR DOWNTO?
				O: OUT STD_LOGIC_VECTOR(0 TO 7));
END DECODER_3_8;

ARCHITECTURE BEHV OF DECODER_3_8 IS
BEGIN
	WITH I SELECT O <=
		"10000000" WHEN "000",
		"01000000" WHEN "001",
		"00100000" WHEN "010",
		"00010000" WHEN "011",
		"00001000" WHEN "100",
		"00000100" WHEN "101",
		"00000010" WHEN "110",
		"00000001" WHEN "111",
		"00000000" WHEN OTHERS;
END BEHV;