LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY ADDER IS
	PORT (X: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
				Y: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
				Z: OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
END ADDER;

ARCHITECTURE BEHV OF ADDER IS
BEGIN
	PROCESS (X,Y)
    VARIABLE C: STD_LOGIC;
  BEGIN
    C := '0';
		FOR I IN 0 TO 15 LOOP
      Z(I) <= X(I) XOR Y(I) XOR C;
      C := (X(I) AND Y(I)) OR (X(I) AND C) OR (Y(I) AND C);
    END LOOP;
  END PROCESS;
END BEHV;