LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY REGISTER_16 IS
	PORT (CLK: IN STD_LOGIC;
	      EN: IN STD_LOGIC;
        D: IN STD_LOGIC_VECTOR(15 downto 0);
        Q: OUT STD_LOGIC_VECTOR(15 downto 0));
END REGISTER_16;

ARCHITECTURE BEHV OF REGISTER_16 IS
BEGIN
	PROCESS (D, CLK, EN)
  BEGIN
    IF EN='1' AND CLK' EVENT AND (NOT (NOT CLK))='1' THEN
			Q <= D;
    END IF;
	END PROCESS;
END BEHV;