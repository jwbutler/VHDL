LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SUB IS
	PORT (X: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
				Y: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
				Z: OUT STD_LOGIC_VECTOR (15 DOWNTO 0));
END SUB;

ARCHITECTURE BEHV OF SUB IS
	BEGIN
	PROCESS (X,Y)
    VARIABLE B: STD_LOGIC;
    BEGIN
	    B := '0';
		FOR I IN 0 TO 15 LOOP
      Z(I) <= X(I) XOR (NOT Y(I)) XOR (NOT B);
			B := (NOT X(I) AND Y(I)) OR (NOT X(I) AND B) OR (Y(I) AND B);
    END LOOP;
  END PROCESS;
END BEHV;